library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity free_run_bin_counter is
	generic (N : integer := 8);
	port (
		clk : in std_logic;
		reset : in std_logic;
		inc, dec : in std_logic;
		enable : in std_logic;
		q : out std_logic_vector(N - 1 downto 0)
	);
end free_run_bin_counter;

architecture arch of free_run_bin_counter is
	signal r_reg : unsigned(N - 1 downto 0);
	signal r_next : unsigned(N - 1 downto 0);
begin
	-- register
	process (clk, reset)
	begin
		if (reset = '1') then
			r_reg <= (others => '0');
		elsif (clk'EVENT and clk = '1') then
			r_reg <= r_next;
		end if;
	end process;
	-- next-state logic
	if inc = '1' then
		r_next <= r_reg + 1;
	elsif dec = '1' then
		r_next <= r_reg - 1;
	else
		r_next <= r_reg;
	end if;
	-- output logic
	q <= std_logic_vector(r_reg);
end arch;